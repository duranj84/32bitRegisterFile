module mux_tb();
	reg [31:0] x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31;
	reg [4:0] select;
	wire [31:0] out;
	
	//COA_Lab3Mux dut (out, x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, select);
	Mux_32x1 dut (x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31, select, out);
	
	initial begin
		select[4:0] <= 5'b00000;
		x0 [31:0] <= 32'd0;
		x1 [31:0] <= 32'd10;
		x2 [31:0] <= 32'd20;
		x3 [31:0] <= 32'd30;
		x4 [31:0] <= 32'd40;
		x5 [31:0] <= 32'd50;
		x6 [31:0] <= 32'd60;
		x7 [31:0] <= 32'd70;
		x8 [31:0] <= 32'd80;
		x9 [31:0] <= 32'd90;
		x10 [31:0] <= 32'd100;
		x11 [31:0] <= 32'd110;
		x12 [31:0] <= 32'd120;
		x13 [31:0] <= 32'd130;
		x14 [31:0] <= 32'd140;
		x15 [31:0] <= 32'd150;
		x16 [31:0] <= 32'd160;
		x17 [31:0] <= 32'd170;
		x18 [31:0] <= 32'd180;
		x19 [31:0] <= 32'd190;
		x20 [31:0] <= 32'd200;
		x21 [31:0] <= 32'd210;
		x22 [31:0] <= 32'd220;
		x23 [31:0] <= 32'd230;
		x24 [31:0] <= 32'd240;
		x25 [31:0] <= 32'd250;
		x26 [31:0] <= 32'd260;
		x27 [31:0] <= 32'd270;
		x28 [31:0] <= 32'd280;
		x29 [31:0] <= 32'd290;
		x30 [31:0] <= 32'd300;
		x31 [31:0] <= 32'd310;
		
	end
	
	always
		#10 select <= select + 1'b1;
		
	initial
		#1000 $stop;

endmodule